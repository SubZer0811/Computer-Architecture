`include "FP_adder.v"

module FP_adder_tb;
reg [31:0]a, b;
wire [31:0]out;
reg clk;

FP_adder FP1 (out, a, b, clk);

initial
begin

	// +ve +ve 
	a = 32'b0_10000000_11110000000000000000000;		// 3.875
	b = 32'b0_10000000_11000000000000000000000;		// 3.5
	// ==> 32'b0_10000001_11011000000000000000000  ans = 7.375

	
	// a = 32'b1_10000000_11100000000000000000000;		// -3.75
	// b = 32'b0_10000000_11000000000000000000000;		// 3.5 // ans:1 01111101 00000000000000000000000
	// // #5 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
	
	
	// // -ve -ve
	// #10 a =	32'b1_10000010_00111000000000000000000;
	// #10 b =	32'b1_10000010_00111000000000000000000;
	// #10 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);

	// #15 a = 32'b0_10000010_00111000000000000000000;
	// #15 b = 32'b0_10000000_11000000000000000000000;
	
	// // infinity case
	//  a = 32'b0_11111111_00000000000000000000000;
	//  b = 32'b1_11111100_00000000000000000000000;

	// #35 a = 32'b0_11111111_00000000000000000000000;
	// #35 b = 32'b0_11111111_00000000000000000000000;

	// #45 a = 32'b0_01111110_01100000000000000000000;
	// #45 b = 32'b1_01111110_00100000000000000000000;
	// // ans:0 01111100 00000000000000000000000

	// // b = 32'b0_01111111_00000000000000000000000;
	// #5 a = 32'h0000;
	// #5 b = 32'h0000;

	#200	$finish();

end

initial begin
	clk = 0;
	forever begin
		#1 clk = ~clk;
	end
end

initial begin
	$monitor("%d# a=%b; b=%b; out=%b", $time, a, b, out);
end

endmodule